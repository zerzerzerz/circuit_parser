module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire net13;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net12;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire net11;
 wire _167_;
 wire _168_;
 wire net10;
 wire net9;
 wire net8;
 wire _172_;
 wire net7;
 wire _174_;
 wire net6;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire net5;
 wire _190_;
 wire _191_;
 wire net4;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire net3;
 wire net2;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire net1;
 wire _235_;
 wire _236_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net54;
 wire net55;
 wire net56;

 INV_X2 _345_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_036_));
 TAPCELL_X1 PHY_14 ();
 NAND2_X1 _347_ (.A1(_036_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_038_));
 INV_X1 _348_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_039_));
 NOR2_X1 _349_ (.A1(_039_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_040_));
 NOR2_X1 _350_ (.A1(_036_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_041_));
 OAI21_X2 _351_ (.A(_038_),
    .B1(_040_),
    .B2(_041_),
    .ZN(_042_));
 INV_X1 _352_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_043_));
 NAND2_X1 _353_ (.A1(_043_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_044_));
 INV_X1 _354_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_045_));
 NAND2_X1 _355_ (.A1(_045_),
    .A2(\dpath.a_lt_b$in1[3] ),
    .ZN(_046_));
 NAND2_X1 _356_ (.A1(_044_),
    .A2(_046_),
    .ZN(_047_));
 INV_X2 _357_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_048_));
 NAND2_X1 _358_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_049_));
 INV_X1 _359_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_050_));
 NAND2_X1 _360_ (.A1(_050_),
    .A2(\dpath.a_lt_b$in1[2] ),
    .ZN(_051_));
 NAND2_X1 _361_ (.A1(_049_),
    .A2(_051_),
    .ZN(_052_));
 NOR2_X1 _362_ (.A1(_047_),
    .A2(_052_),
    .ZN(_053_));
 NAND2_X1 _363_ (.A1(_042_),
    .A2(_053_),
    .ZN(_054_));
 INV_X1 _364_ (.A(_046_),
    .ZN(_055_));
 OAI21_X1 _365_ (.A(_044_),
    .B1(_055_),
    .B2(_049_),
    .ZN(_056_));
 INV_X1 _366_ (.A(_056_),
    .ZN(_057_));
 NAND2_X2 _367_ (.A1(_054_),
    .A2(_057_),
    .ZN(_058_));
 TAPCELL_X1 PHY_13 ();
 XNOR2_X1 _369_ (.A(\dpath.a_lt_b$in1[5] ),
    .B(\dpath.a_lt_b$in0[5] ),
    .ZN(_060_));
 XNOR2_X2 _370_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .ZN(_061_));
 NAND2_X1 _371_ (.A1(_060_),
    .A2(_061_),
    .ZN(_062_));
 XNOR2_X1 _372_ (.A(\dpath.a_lt_b$in1[7] ),
    .B(\dpath.a_lt_b$in0[7] ),
    .ZN(_063_));
 XNOR2_X2 _373_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .ZN(_064_));
 NAND2_X4 _374_ (.A1(_063_),
    .A2(_064_),
    .ZN(_065_));
 NOR2_X4 _375_ (.A1(_062_),
    .A2(_065_),
    .ZN(_066_));
 NAND2_X4 _376_ (.A1(_058_),
    .A2(_066_),
    .ZN(_067_));
 INV_X1 _377_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_068_));
 NAND2_X1 _378_ (.A1(_068_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_069_));
 INV_X1 _379_ (.A(\dpath.a_lt_b$in0[5] ),
    .ZN(_070_));
 OAI21_X1 _380_ (.A(_069_),
    .B1(\dpath.a_lt_b$in1[5] ),
    .B2(_070_),
    .ZN(_071_));
 INV_X1 _381_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_072_));
 NOR2_X1 _382_ (.A1(_072_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_073_));
 INV_X1 _383_ (.A(_073_),
    .ZN(_074_));
 NAND2_X1 _384_ (.A1(_071_),
    .A2(_074_),
    .ZN(_075_));
 NOR2_X4 _385_ (.A1(_075_),
    .A2(_065_),
    .ZN(_076_));
 INV_X1 _386_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_077_));
 NAND2_X1 _387_ (.A1(_077_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_078_));
 INV_X2 _388_ (.A(_063_),
    .ZN(_079_));
 INV_X1 _389_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_080_));
 NAND2_X1 _390_ (.A1(_080_),
    .A2(net56),
    .ZN(_081_));
 OAI21_X1 _391_ (.A(_078_),
    .B1(_079_),
    .B2(_081_),
    .ZN(_082_));
 NOR2_X2 _392_ (.A1(_076_),
    .A2(_082_),
    .ZN(_083_));
 NAND2_X4 _393_ (.A1(_067_),
    .A2(_083_),
    .ZN(_084_));
 INV_X2 _394_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_085_));
 XNOR2_X2 _395_ (.A(_085_),
    .B(\dpath.a_lt_b$in0[11] ),
    .ZN(_086_));
 INV_X2 _396_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_087_));
 XNOR2_X1 _397_ (.A(_087_),
    .B(\dpath.a_lt_b$in0[10] ),
    .ZN(_088_));
 NOR2_X1 _398_ (.A1(_086_),
    .A2(_088_),
    .ZN(_089_));
 XNOR2_X2 _399_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .ZN(_090_));
 XNOR2_X2 _400_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in0[8] ),
    .ZN(_091_));
 NAND2_X1 _401_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 INV_X1 _402_ (.A(_092_),
    .ZN(_093_));
 AND2_X1 _403_ (.A1(_089_),
    .A2(_093_),
    .ZN(_094_));
 NAND2_X4 _404_ (.A1(_084_),
    .A2(_094_),
    .ZN(_095_));
 NAND2_X1 _405_ (.A1(_085_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_096_));
 NAND2_X1 _406_ (.A1(_087_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_097_));
 OAI21_X1 _407_ (.A(_096_),
    .B1(_086_),
    .B2(_097_),
    .ZN(_098_));
 INV_X1 _408_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_099_));
 NOR2_X1 _409_ (.A1(_099_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_100_));
 INV_X1 _410_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_101_));
 AND2_X1 _411_ (.A1(_101_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_102_));
 AOI21_X1 _412_ (.A(_100_),
    .B1(_090_),
    .B2(_102_),
    .ZN(_103_));
 INV_X1 _413_ (.A(_103_),
    .ZN(_104_));
 AOI21_X2 _414_ (.A(_098_),
    .B1(_104_),
    .B2(_089_),
    .ZN(_105_));
 NAND2_X4 _415_ (.A1(_095_),
    .A2(_105_),
    .ZN(_106_));
 XNOR2_X2 _416_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in0[12] ),
    .ZN(_107_));
 INV_X1 _417_ (.A(_107_),
    .ZN(_108_));
 INV_X2 _418_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_109_));
 XNOR2_X2 _419_ (.A(_109_),
    .B(\dpath.a_lt_b$in0[13] ),
    .ZN(_110_));
 NOR2_X1 _420_ (.A1(_108_),
    .A2(_110_),
    .ZN(_111_));
 NAND2_X4 _421_ (.A1(_106_),
    .A2(_111_),
    .ZN(_112_));
 NAND2_X1 _422_ (.A1(_109_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_113_));
 INV_X1 _423_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_114_));
 NAND2_X1 _424_ (.A1(_114_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_115_));
 OAI21_X1 _425_ (.A(_113_),
    .B1(_110_),
    .B2(_115_),
    .ZN(_116_));
 INV_X1 _426_ (.A(_116_),
    .ZN(_117_));
 NAND2_X4 _427_ (.A1(_112_),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _428_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_119_));
 XNOR2_X1 _429_ (.A(_119_),
    .B(\dpath.a_lt_b$in0[14] ),
    .ZN(_120_));
 INV_X1 _430_ (.A(_120_),
    .ZN(_121_));
 NAND2_X4 _431_ (.A1(_118_),
    .A2(_121_),
    .ZN(_122_));
 NAND2_X1 _432_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_123_));
 NAND2_X4 _433_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 INV_X2 _434_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_125_));
 XNOR2_X2 _435_ (.A(_125_),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_126_));
 INV_X1 _436_ (.A(_126_),
    .ZN(_127_));
 NAND2_X4 _437_ (.A1(_124_),
    .A2(_127_),
    .ZN(_128_));
 NAND3_X2 _438_ (.A1(_122_),
    .A2(_123_),
    .A3(_126_),
    .ZN(_129_));
 AND2_X4 _439_ (.A1(_128_),
    .A2(_129_),
    .ZN(net43));
 XNOR2_X1 _440_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .ZN(_130_));
 INV_X1 _441_ (.A(_040_),
    .ZN(_131_));
 XNOR2_X1 _442_ (.A(_130_),
    .B(_131_),
    .ZN(_132_));
 INV_X1 _443_ (.A(_132_),
    .ZN(net44));
 INV_X1 _444_ (.A(_052_),
    .ZN(_133_));
 XNOR2_X1 _445_ (.A(_042_),
    .B(_133_),
    .ZN(_134_));
 INV_X1 _446_ (.A(_134_),
    .ZN(net45));
 NAND2_X1 _447_ (.A1(_042_),
    .A2(_133_),
    .ZN(_135_));
 NAND2_X1 _448_ (.A1(_135_),
    .A2(_049_),
    .ZN(_136_));
 XNOR2_X1 _449_ (.A(_136_),
    .B(_047_),
    .ZN(net46));
 XNOR2_X1 _450_ (.A(_058_),
    .B(_061_),
    .ZN(_137_));
 INV_X1 _451_ (.A(_137_),
    .ZN(net47));
 NAND2_X1 _452_ (.A1(_058_),
    .A2(_061_),
    .ZN(_138_));
 NAND2_X1 _453_ (.A1(_138_),
    .A2(_069_),
    .ZN(_139_));
 XOR2_X1 _454_ (.A(_139_),
    .B(_060_),
    .Z(net48));
 INV_X1 _455_ (.A(_071_),
    .ZN(_140_));
 AOI21_X1 _456_ (.A(_073_),
    .B1(_138_),
    .B2(_140_),
    .ZN(_141_));
 XNOR2_X1 _457_ (.A(_141_),
    .B(_064_),
    .ZN(_142_));
 INV_X1 _458_ (.A(_142_),
    .ZN(net49));
 NAND2_X1 _459_ (.A1(_141_),
    .A2(_064_),
    .ZN(_143_));
 NAND2_X1 _460_ (.A1(_143_),
    .A2(_081_),
    .ZN(_144_));
 XNOR2_X1 _461_ (.A(_144_),
    .B(_079_),
    .ZN(net50));
 XNOR2_X1 _462_ (.A(_084_),
    .B(_091_),
    .ZN(_145_));
 INV_X1 _463_ (.A(_145_),
    .ZN(net51));
 AOI21_X1 _464_ (.A(_102_),
    .B1(_084_),
    .B2(_091_),
    .ZN(_146_));
 XNOR2_X1 _465_ (.A(_146_),
    .B(_090_),
    .ZN(net52));
 NAND2_X1 _466_ (.A1(_084_),
    .A2(_093_),
    .ZN(_147_));
 NAND2_X1 _467_ (.A1(_147_),
    .A2(_103_),
    .ZN(_148_));
 INV_X1 _468_ (.A(_088_),
    .ZN(_149_));
 XNOR2_X1 _469_ (.A(_148_),
    .B(_149_),
    .ZN(_150_));
 INV_X1 _470_ (.A(_150_),
    .ZN(net38));
 NAND2_X1 _471_ (.A1(_148_),
    .A2(_149_),
    .ZN(_151_));
 NAND2_X1 _472_ (.A1(_151_),
    .A2(_097_),
    .ZN(_152_));
 XNOR2_X1 _473_ (.A(_152_),
    .B(_086_),
    .ZN(net39));
 XNOR2_X1 _474_ (.A(_106_),
    .B(_107_),
    .ZN(_153_));
 INV_X1 _475_ (.A(_153_),
    .ZN(net40));
 NAND2_X1 _476_ (.A1(_106_),
    .A2(_107_),
    .ZN(_154_));
 NAND2_X1 _477_ (.A1(_154_),
    .A2(_115_),
    .ZN(_155_));
 XNOR2_X1 _478_ (.A(_155_),
    .B(_110_),
    .ZN(net41));
 XNOR2_X1 _479_ (.A(_118_),
    .B(_121_),
    .ZN(_156_));
 INV_X1 _480_ (.A(_156_),
    .ZN(net42));
 XNOR2_X1 _481_ (.A(_039_),
    .B(\dpath.a_lt_b$in0[0] ),
    .ZN(net37));
 NAND4_X1 _482_ (.A1(_119_),
    .A2(_125_),
    .A3(_039_),
    .A4(_036_),
    .ZN(_157_));
 NAND3_X1 _483_ (.A1(_087_),
    .A2(_085_),
    .A3(_114_),
    .ZN(_158_));
 NOR3_X1 _484_ (.A1(_157_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .A3(_158_),
    .ZN(_159_));
 INV_X1 _485_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_160_));
 NAND4_X1 _486_ (.A1(_080_),
    .A2(_077_),
    .A3(_101_),
    .A4(_160_),
    .ZN(_161_));
 NAND4_X1 _487_ (.A1(_048_),
    .A2(_043_),
    .A3(_068_),
    .A4(_072_),
    .ZN(_162_));
 NOR2_X1 _488_ (.A1(_161_),
    .A2(_162_),
    .ZN(_163_));
 NAND2_X1 _489_ (.A1(_159_),
    .A2(_163_),
    .ZN(_164_));
 INV_X1 _490_ (.A(_164_),
    .ZN(_165_));
 TAPCELL_X1 PHY_12 ();
 INV_X1 _492_ (.A(\ctrl.state.out[2] ),
    .ZN(_167_));
 OR2_X1 _493_ (.A1(_167_),
    .A2(net34),
    .ZN(_168_));
 TAPCELL_X1 PHY_11 ();
 TAPCELL_X1 PHY_10 ();
 TAPCELL_X1 PHY_9 ();
 NAND2_X1 _497_ (.A1(net36),
    .A2(net33),
    .ZN(_172_));
 OAI22_X1 _498_ (.A1(_165_),
    .A2(_168_),
    .B1(net34),
    .B2(_172_),
    .ZN(_002_));
 TAPCELL_X1 PHY_8 ();
 AND3_X1 _500_ (.A1(_167_),
    .A2(_003_),
    .A3(\ctrl.state.out[1] ),
    .ZN(net53));
 AOI21_X1 _501_ (.A(net34),
    .B1(net53),
    .B2(net35),
    .ZN(_174_));
 TAPCELL_X1 PHY_7 ();
 INV_X1 _503_ (.A(net36),
    .ZN(_176_));
 OAI21_X1 _504_ (.A(_174_),
    .B1(_176_),
    .B2(net33),
    .ZN(_000_));
 NAND2_X1 _505_ (.A1(_174_),
    .A2(\ctrl.state.out[1] ),
    .ZN(_177_));
 OAI21_X1 _506_ (.A(_177_),
    .B1(_164_),
    .B2(_168_),
    .ZN(_001_));
 NAND2_X1 _507_ (.A1(_125_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_178_));
 OAI21_X1 _508_ (.A(_178_),
    .B1(_126_),
    .B2(_123_),
    .ZN(_179_));
 NOR2_X1 _509_ (.A1(_120_),
    .A2(_126_),
    .ZN(_180_));
 AOI21_X1 _510_ (.A(_179_),
    .B1(_116_),
    .B2(_180_),
    .ZN(_181_));
 NAND2_X1 _511_ (.A1(_111_),
    .A2(_180_),
    .ZN(_182_));
 OAI21_X1 _512_ (.A(_181_),
    .B1(_105_),
    .B2(_182_),
    .ZN(_183_));
 INV_X2 _513_ (.A(_183_),
    .ZN(_184_));
 INV_X1 _514_ (.A(_182_),
    .ZN(_185_));
 NAND3_X2 _515_ (.A1(_084_),
    .A2(_094_),
    .A3(_185_),
    .ZN(_186_));
 NAND3_X1 _516_ (.A1(_184_),
    .A2(_186_),
    .A3(\ctrl.state.out[2] ),
    .ZN(_187_));
 NAND2_X4 _517_ (.A1(_187_),
    .A2(_003_),
    .ZN(_188_));
 TAPCELL_X1 PHY_6 ();
 MUX2_X1 _519_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(net1),
    .S(net36),
    .Z(_190_));
 NAND2_X1 _520_ (.A1(_188_),
    .A2(_190_),
    .ZN(_191_));
 TAPCELL_X1 PHY_5 ();
 OAI21_X1 _522_ (.A(_191_),
    .B1(_039_),
    .B2(_188_),
    .ZN(_004_));
 MUX2_X1 _523_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(net12),
    .S(net36),
    .Z(_193_));
 NAND2_X1 _524_ (.A1(_188_),
    .A2(_193_),
    .ZN(_194_));
 OAI21_X1 _525_ (.A(_194_),
    .B1(_036_),
    .B2(_188_),
    .ZN(_005_));
 NAND2_X1 _526_ (.A1(net36),
    .A2(net23),
    .ZN(_195_));
 OAI21_X1 _527_ (.A(_195_),
    .B1(net36),
    .B2(_050_),
    .ZN(_196_));
 NAND2_X1 _528_ (.A1(_188_),
    .A2(_196_),
    .ZN(_197_));
 OAI21_X1 _529_ (.A(_197_),
    .B1(_048_),
    .B2(_188_),
    .ZN(_006_));
 NAND2_X1 _530_ (.A1(net36),
    .A2(net26),
    .ZN(_198_));
 OAI21_X1 _531_ (.A(_198_),
    .B1(net36),
    .B2(_045_),
    .ZN(_199_));
 NAND2_X1 _532_ (.A1(_188_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _533_ (.A(_200_),
    .B1(_043_),
    .B2(_188_),
    .ZN(_007_));
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_3 ();
 MUX2_X1 _536_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(net27),
    .S(net36),
    .Z(_203_));
 NAND2_X1 _537_ (.A1(_188_),
    .A2(_203_),
    .ZN(_204_));
 OAI21_X1 _538_ (.A(_204_),
    .B1(_068_),
    .B2(_188_),
    .ZN(_008_));
 NAND2_X1 _539_ (.A1(net36),
    .A2(net28),
    .ZN(_205_));
 OAI21_X1 _540_ (.A(_205_),
    .B1(net36),
    .B2(_070_),
    .ZN(_206_));
 NAND2_X1 _541_ (.A1(_188_),
    .A2(_206_),
    .ZN(_207_));
 OAI21_X1 _542_ (.A(_207_),
    .B1(_072_),
    .B2(_188_),
    .ZN(_009_));
 MUX2_X1 _543_ (.A(net55),
    .B(net29),
    .S(net36),
    .Z(_208_));
 NAND2_X1 _544_ (.A1(_188_),
    .A2(_208_),
    .ZN(_209_));
 OAI21_X1 _545_ (.A(_209_),
    .B1(_080_),
    .B2(_188_),
    .ZN(_010_));
 MUX2_X1 _546_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(net30),
    .S(net36),
    .Z(_210_));
 NAND2_X1 _547_ (.A1(_188_),
    .A2(_210_),
    .ZN(_211_));
 OAI21_X1 _548_ (.A(_211_),
    .B1(_077_),
    .B2(_188_),
    .ZN(_011_));
 MUX2_X1 _549_ (.A(\dpath.a_lt_b$in0[8] ),
    .B(net31),
    .S(net36),
    .Z(_212_));
 NAND2_X1 _550_ (.A1(_188_),
    .A2(_212_),
    .ZN(_213_));
 OAI21_X1 _551_ (.A(_213_),
    .B1(_101_),
    .B2(_188_),
    .ZN(_012_));
 NAND2_X1 _552_ (.A1(net36),
    .A2(net32),
    .ZN(_214_));
 OAI21_X1 _553_ (.A(_214_),
    .B1(net36),
    .B2(_099_),
    .ZN(_215_));
 NAND2_X1 _554_ (.A1(_188_),
    .A2(_215_),
    .ZN(_216_));
 OAI21_X1 _555_ (.A(_216_),
    .B1(_160_),
    .B2(_188_),
    .ZN(_013_));
 MUX2_X1 _556_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(net2),
    .S(net36),
    .Z(_217_));
 NAND2_X1 _557_ (.A1(_188_),
    .A2(_217_),
    .ZN(_218_));
 OAI21_X1 _558_ (.A(_218_),
    .B1(_087_),
    .B2(_188_),
    .ZN(_014_));
 MUX2_X1 _559_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(net3),
    .S(net36),
    .Z(_219_));
 NAND2_X1 _560_ (.A1(_188_),
    .A2(_219_),
    .ZN(_220_));
 OAI21_X1 _561_ (.A(_220_),
    .B1(_085_),
    .B2(_188_),
    .ZN(_015_));
 MUX2_X1 _562_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(net4),
    .S(net36),
    .Z(_221_));
 NAND2_X1 _563_ (.A1(_188_),
    .A2(_221_),
    .ZN(_222_));
 OAI21_X1 _564_ (.A(_222_),
    .B1(_114_),
    .B2(_188_),
    .ZN(_016_));
 MUX2_X1 _565_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(net5),
    .S(net36),
    .Z(_223_));
 NAND2_X1 _566_ (.A1(_188_),
    .A2(_223_),
    .ZN(_224_));
 OAI21_X1 _567_ (.A(_224_),
    .B1(_109_),
    .B2(_188_),
    .ZN(_017_));
 MUX2_X1 _568_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(net6),
    .S(net36),
    .Z(_225_));
 NAND2_X1 _569_ (.A1(_188_),
    .A2(_225_),
    .ZN(_226_));
 OAI21_X1 _570_ (.A(_226_),
    .B1(_119_),
    .B2(_188_),
    .ZN(_018_));
 MUX2_X1 _571_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(net7),
    .S(net36),
    .Z(_227_));
 NAND2_X1 _572_ (.A1(_188_),
    .A2(_227_),
    .ZN(_228_));
 OAI21_X1 _573_ (.A(_228_),
    .B1(_125_),
    .B2(_188_),
    .ZN(_019_));
 NAND2_X1 _574_ (.A1(_184_),
    .A2(_186_),
    .ZN(_229_));
 NAND3_X4 _575_ (.A1(_229_),
    .A2(\ctrl.state.out[2] ),
    .A3(_003_),
    .ZN(_230_));
 INV_X8 _576_ (.A(_230_),
    .ZN(_231_));
 NAND2_X1 _577_ (.A1(_231_),
    .A2(net37),
    .ZN(_232_));
 NAND4_X4 _578_ (.A1(_184_),
    .A2(_186_),
    .A3(\ctrl.state.out[2] ),
    .A4(_003_),
    .ZN(_233_));
 TAPCELL_X1 PHY_2 ();
 OAI21_X1 _580_ (.A(_232_),
    .B1(_233_),
    .B2(_039_),
    .ZN(_235_));
 NOR2_X4 _581_ (.A1(_167_),
    .A2(net36),
    .ZN(_236_));
 TAPCELL_X1 PHY_1 ();
 NAND2_X1 _583_ (.A1(_235_),
    .A2(_236_),
    .ZN(_238_));
 NAND2_X1 _584_ (.A1(net36),
    .A2(net8),
    .ZN(_239_));
 NOR2_X4 _585_ (.A1(\ctrl.state.out[2] ),
    .A2(net36),
    .ZN(_240_));
 TAPCELL_X1 PHY_0 ();
 NAND2_X1 _587_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_242_));
 NAND3_X1 _588_ (.A1(_238_),
    .A2(_239_),
    .A3(_242_),
    .ZN(_020_));
 OAI22_X1 _589_ (.A1(_233_),
    .A2(_036_),
    .B1(_230_),
    .B2(_132_),
    .ZN(_243_));
 NAND2_X1 _590_ (.A1(_243_),
    .A2(_236_),
    .ZN(_244_));
 NAND2_X1 _591_ (.A1(net36),
    .A2(net9),
    .ZN(_245_));
 NAND2_X1 _592_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_246_));
 NAND3_X1 _593_ (.A1(_244_),
    .A2(_245_),
    .A3(_246_),
    .ZN(_021_));
 OAI22_X1 _594_ (.A1(_233_),
    .A2(_048_),
    .B1(_230_),
    .B2(_134_),
    .ZN(_247_));
 NAND2_X1 _595_ (.A1(_247_),
    .A2(_236_),
    .ZN(_248_));
 NAND2_X1 _596_ (.A1(net10),
    .A2(net36),
    .ZN(_249_));
 NAND2_X1 _597_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_250_));
 NAND3_X1 _598_ (.A1(_248_),
    .A2(_249_),
    .A3(_250_),
    .ZN(_022_));
 NAND2_X1 _599_ (.A1(_231_),
    .A2(net46),
    .ZN(_251_));
 OAI21_X1 _600_ (.A(_251_),
    .B1(_233_),
    .B2(_043_),
    .ZN(_252_));
 NAND2_X1 _601_ (.A1(_252_),
    .A2(_236_),
    .ZN(_253_));
 NAND2_X1 _602_ (.A1(net11),
    .A2(net36),
    .ZN(_254_));
 NAND2_X1 _603_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_255_));
 NAND3_X1 _604_ (.A1(_253_),
    .A2(_254_),
    .A3(_255_),
    .ZN(_023_));
 OAI22_X1 _605_ (.A1(_233_),
    .A2(_068_),
    .B1(_230_),
    .B2(_137_),
    .ZN(_256_));
 NAND2_X1 _606_ (.A1(_256_),
    .A2(_236_),
    .ZN(_257_));
 NAND2_X1 _607_ (.A1(net13),
    .A2(net36),
    .ZN(_258_));
 NAND2_X1 _608_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_259_));
 NAND3_X1 _609_ (.A1(_257_),
    .A2(_258_),
    .A3(_259_),
    .ZN(_024_));
 NAND2_X1 _610_ (.A1(_231_),
    .A2(net48),
    .ZN(_260_));
 OAI21_X1 _611_ (.A(_260_),
    .B1(_233_),
    .B2(_072_),
    .ZN(_261_));
 NAND2_X1 _612_ (.A1(_261_),
    .A2(_236_),
    .ZN(_262_));
 NAND2_X1 _613_ (.A1(net14),
    .A2(net36),
    .ZN(_263_));
 NAND2_X1 _614_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_264_));
 NAND3_X1 _615_ (.A1(_262_),
    .A2(_263_),
    .A3(_264_),
    .ZN(_025_));
 OAI22_X1 _616_ (.A1(_233_),
    .A2(_080_),
    .B1(_230_),
    .B2(_142_),
    .ZN(_265_));
 NAND2_X1 _617_ (.A1(_265_),
    .A2(_236_),
    .ZN(_266_));
 NAND2_X1 _618_ (.A1(net15),
    .A2(net36),
    .ZN(_267_));
 NAND2_X1 _619_ (.A1(_240_),
    .A2(net54),
    .ZN(_268_));
 NAND3_X1 _620_ (.A1(_266_),
    .A2(_267_),
    .A3(_268_),
    .ZN(_026_));
 NAND2_X1 _621_ (.A1(net50),
    .A2(_231_),
    .ZN(_269_));
 OAI21_X1 _622_ (.A(_269_),
    .B1(_077_),
    .B2(_233_),
    .ZN(_270_));
 NAND2_X1 _623_ (.A1(_270_),
    .A2(_236_),
    .ZN(_271_));
 NAND2_X1 _624_ (.A1(net16),
    .A2(net36),
    .ZN(_272_));
 NAND2_X1 _625_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_273_));
 NAND3_X1 _626_ (.A1(_271_),
    .A2(_272_),
    .A3(_273_),
    .ZN(_027_));
 OAI22_X1 _627_ (.A1(_233_),
    .A2(_101_),
    .B1(_230_),
    .B2(_145_),
    .ZN(_274_));
 NAND2_X1 _628_ (.A1(_274_),
    .A2(_236_),
    .ZN(_275_));
 NAND2_X1 _629_ (.A1(net17),
    .A2(net36),
    .ZN(_276_));
 NAND2_X1 _630_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_277_));
 NAND3_X1 _631_ (.A1(_275_),
    .A2(_276_),
    .A3(_277_),
    .ZN(_028_));
 NAND2_X1 _632_ (.A1(_231_),
    .A2(net52),
    .ZN(_278_));
 OAI21_X1 _633_ (.A(_278_),
    .B1(_233_),
    .B2(_160_),
    .ZN(_279_));
 NAND2_X1 _634_ (.A1(_279_),
    .A2(_236_),
    .ZN(_280_));
 NAND2_X1 _635_ (.A1(net18),
    .A2(net36),
    .ZN(_281_));
 NAND2_X1 _636_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_282_));
 NAND3_X1 _637_ (.A1(_280_),
    .A2(_281_),
    .A3(_282_),
    .ZN(_029_));
 OAI22_X1 _638_ (.A1(_150_),
    .A2(_230_),
    .B1(_233_),
    .B2(_087_),
    .ZN(_283_));
 NAND2_X1 _639_ (.A1(_283_),
    .A2(_236_),
    .ZN(_284_));
 NAND2_X1 _640_ (.A1(net19),
    .A2(net36),
    .ZN(_285_));
 NAND2_X1 _641_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_286_));
 NAND3_X1 _642_ (.A1(_284_),
    .A2(_285_),
    .A3(_286_),
    .ZN(_030_));
 NAND2_X1 _643_ (.A1(net39),
    .A2(_231_),
    .ZN(_287_));
 OAI21_X1 _644_ (.A(_287_),
    .B1(_085_),
    .B2(_233_),
    .ZN(_288_));
 NAND2_X1 _645_ (.A1(_288_),
    .A2(_236_),
    .ZN(_289_));
 AND2_X1 _646_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_290_));
 AOI21_X1 _647_ (.A(_290_),
    .B1(net20),
    .B2(net36),
    .ZN(_291_));
 NAND2_X1 _648_ (.A1(_289_),
    .A2(_291_),
    .ZN(_031_));
 OAI22_X1 _649_ (.A1(_153_),
    .A2(_230_),
    .B1(_233_),
    .B2(_114_),
    .ZN(_292_));
 NAND2_X1 _650_ (.A1(_292_),
    .A2(_236_),
    .ZN(_293_));
 NAND2_X1 _651_ (.A1(net21),
    .A2(net36),
    .ZN(_294_));
 NAND2_X1 _652_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_295_));
 NAND3_X1 _653_ (.A1(_293_),
    .A2(_294_),
    .A3(_295_),
    .ZN(_032_));
 NAND2_X1 _654_ (.A1(net41),
    .A2(_231_),
    .ZN(_296_));
 OAI21_X1 _655_ (.A(_296_),
    .B1(_109_),
    .B2(_233_),
    .ZN(_297_));
 NAND2_X1 _656_ (.A1(_297_),
    .A2(_236_),
    .ZN(_298_));
 AND2_X1 _657_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_299_));
 AOI21_X1 _658_ (.A(_299_),
    .B1(net22),
    .B2(net36),
    .ZN(_300_));
 NAND2_X1 _659_ (.A1(_298_),
    .A2(_300_),
    .ZN(_033_));
 OAI22_X1 _660_ (.A1(_156_),
    .A2(_230_),
    .B1(_233_),
    .B2(_119_),
    .ZN(_301_));
 NAND2_X1 _661_ (.A1(_301_),
    .A2(_236_),
    .ZN(_302_));
 AND2_X1 _662_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_303_));
 AOI21_X1 _663_ (.A(_303_),
    .B1(net24),
    .B2(net36),
    .ZN(_304_));
 NAND2_X1 _664_ (.A1(_302_),
    .A2(_304_),
    .ZN(_034_));
 NAND3_X1 _665_ (.A1(_128_),
    .A2(_129_),
    .A3(_231_),
    .ZN(_305_));
 OR2_X1 _666_ (.A1(_233_),
    .A2(_125_),
    .ZN(_306_));
 NAND2_X1 _667_ (.A1(_305_),
    .A2(_306_),
    .ZN(_307_));
 NAND2_X1 _668_ (.A1(_307_),
    .A2(_236_),
    .ZN(_308_));
 AND2_X1 _669_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_309_));
 AOI21_X1 _670_ (.A(_309_),
    .B1(net25),
    .B2(net36),
    .ZN(_310_));
 NAND2_X1 _671_ (.A1(_308_),
    .A2(_310_),
    .ZN(_035_));
 DFF_X2 _672_ (.D(_000_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net36),
    .QN(_003_));
 DFF_X1 _673_ (.D(_001_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_344_));
 DFF_X2 _674_ (.D(_002_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_343_));
 DFF_X1 _675_ (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_342_));
 DFF_X1 _676_ (.D(_005_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_341_));
 DFF_X1 _677_ (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_340_));
 DFF_X1 _678_ (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_339_));
 DFF_X1 _679_ (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_338_));
 DFF_X1 _680_ (.D(_009_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_337_));
 DFF_X1 _681_ (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_336_));
 DFF_X1 _682_ (.D(_011_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_335_));
 DFF_X1 _683_ (.D(_012_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_334_));
 DFF_X1 _684_ (.D(_013_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_333_));
 DFF_X1 _685_ (.D(_014_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_332_));
 DFF_X1 _686_ (.D(_015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_331_));
 DFF_X1 _687_ (.D(_016_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_330_));
 DFF_X1 _688_ (.D(_017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_329_));
 DFF_X1 _689_ (.D(_018_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_328_));
 DFF_X1 _690_ (.D(_019_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_327_));
 DFF_X1 _691_ (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_326_));
 DFF_X2 _692_ (.D(_021_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_325_));
 DFF_X1 _693_ (.D(_022_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_324_));
 DFF_X1 _694_ (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_323_));
 DFF_X2 _695_ (.D(_024_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_322_));
 DFF_X1 _696_ (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_321_));
 DFF_X2 _697_ (.D(_026_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_320_));
 DFF_X1 _698_ (.D(_027_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_319_));
 DFF_X2 _699_ (.D(_028_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_318_));
 DFF_X2 _700_ (.D(_029_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_317_));
 DFF_X1 _701_ (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_316_));
 DFF_X2 _702_ (.D(_031_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_315_));
 DFF_X2 _703_ (.D(_032_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_314_));
 DFF_X2 _704_ (.D(_033_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_313_));
 DFF_X1 _705_ (.D(_034_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_312_));
 DFF_X2 _706_ (.D(_035_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_311_));
 TAPCELL_X1 PHY_15 ();
 TAPCELL_X1 PHY_16 ();
 TAPCELL_X1 PHY_17 ();
 TAPCELL_X1 PHY_18 ();
 TAPCELL_X1 PHY_19 ();
 TAPCELL_X1 PHY_20 ();
 TAPCELL_X1 PHY_21 ();
 TAPCELL_X1 PHY_22 ();
 TAPCELL_X1 PHY_23 ();
 TAPCELL_X1 PHY_24 ();
 TAPCELL_X1 PHY_25 ();
 TAPCELL_X1 PHY_26 ();
 TAPCELL_X1 PHY_27 ();
 TAPCELL_X1 PHY_28 ();
 TAPCELL_X1 PHY_29 ();
 TAPCELL_X1 PHY_30 ();
 TAPCELL_X1 PHY_31 ();
 TAPCELL_X1 PHY_32 ();
 TAPCELL_X1 PHY_33 ();
 TAPCELL_X1 PHY_34 ();
 TAPCELL_X1 PHY_35 ();
 TAPCELL_X1 PHY_36 ();
 TAPCELL_X1 PHY_37 ();
 TAPCELL_X1 PHY_38 ();
 TAPCELL_X1 PHY_39 ();
 TAPCELL_X1 PHY_40 ();
 TAPCELL_X1 PHY_41 ();
 TAPCELL_X1 PHY_42 ();
 TAPCELL_X1 PHY_43 ();
 TAPCELL_X1 PHY_44 ();
 TAPCELL_X1 PHY_45 ();
 TAPCELL_X1 PHY_46 ();
 TAPCELL_X1 PHY_47 ();
 TAPCELL_X1 PHY_48 ();
 TAPCELL_X1 PHY_49 ();
 TAPCELL_X1 PHY_50 ();
 TAPCELL_X1 PHY_51 ();
 TAPCELL_X1 PHY_52 ();
 TAPCELL_X1 PHY_53 ();
 TAPCELL_X1 PHY_54 ();
 TAPCELL_X1 PHY_55 ();
 TAPCELL_X1 PHY_56 ();
 TAPCELL_X1 PHY_57 ();
 TAPCELL_X1 PHY_58 ();
 TAPCELL_X1 PHY_59 ();
 TAPCELL_X1 PHY_60 ();
 TAPCELL_X1 PHY_61 ();
 TAPCELL_X1 PHY_62 ();
 TAPCELL_X1 PHY_63 ();
 TAPCELL_X1 PHY_64 ();
 TAPCELL_X1 PHY_65 ();
 TAPCELL_X1 PHY_66 ();
 TAPCELL_X1 PHY_67 ();
 TAPCELL_X1 PHY_68 ();
 TAPCELL_X1 PHY_69 ();
 BUF_X1 input1 (.A(req_msg[0]),
    .Z(net1));
 BUF_X1 input2 (.A(req_msg[10]),
    .Z(net2));
 BUF_X1 input3 (.A(req_msg[11]),
    .Z(net3));
 BUF_X1 input4 (.A(req_msg[12]),
    .Z(net4));
 BUF_X1 input5 (.A(req_msg[13]),
    .Z(net5));
 BUF_X1 input6 (.A(req_msg[14]),
    .Z(net6));
 BUF_X1 input7 (.A(req_msg[15]),
    .Z(net7));
 BUF_X1 input8 (.A(req_msg[16]),
    .Z(net8));
 BUF_X1 input9 (.A(req_msg[17]),
    .Z(net9));
 BUF_X1 input10 (.A(req_msg[18]),
    .Z(net10));
 BUF_X1 input11 (.A(req_msg[19]),
    .Z(net11));
 BUF_X1 input12 (.A(req_msg[1]),
    .Z(net12));
 BUF_X1 input13 (.A(req_msg[20]),
    .Z(net13));
 BUF_X1 input14 (.A(req_msg[21]),
    .Z(net14));
 BUF_X1 input15 (.A(req_msg[22]),
    .Z(net15));
 BUF_X1 input16 (.A(req_msg[23]),
    .Z(net16));
 BUF_X1 input17 (.A(req_msg[24]),
    .Z(net17));
 BUF_X1 input18 (.A(req_msg[25]),
    .Z(net18));
 BUF_X1 input19 (.A(req_msg[26]),
    .Z(net19));
 BUF_X1 input20 (.A(req_msg[27]),
    .Z(net20));
 BUF_X1 input21 (.A(req_msg[28]),
    .Z(net21));
 BUF_X1 input22 (.A(req_msg[29]),
    .Z(net22));
 BUF_X1 input23 (.A(req_msg[2]),
    .Z(net23));
 BUF_X1 input24 (.A(req_msg[30]),
    .Z(net24));
 BUF_X1 input25 (.A(req_msg[31]),
    .Z(net25));
 BUF_X1 input26 (.A(req_msg[3]),
    .Z(net26));
 BUF_X1 input27 (.A(req_msg[4]),
    .Z(net27));
 BUF_X1 input28 (.A(req_msg[5]),
    .Z(net28));
 BUF_X1 input29 (.A(req_msg[6]),
    .Z(net29));
 BUF_X1 input30 (.A(req_msg[7]),
    .Z(net30));
 BUF_X1 input31 (.A(req_msg[8]),
    .Z(net31));
 BUF_X1 input32 (.A(req_msg[9]),
    .Z(net32));
 BUF_X1 input33 (.A(req_val),
    .Z(net33));
 BUF_X1 input34 (.A(reset),
    .Z(net34));
 BUF_X1 input35 (.A(resp_rdy),
    .Z(net35));
 BUF_X1 output36 (.A(net36),
    .Z(req_rdy));
 BUF_X1 output37 (.A(net37),
    .Z(resp_msg[0]));
 BUF_X1 output38 (.A(net38),
    .Z(resp_msg[10]));
 BUF_X1 output39 (.A(net39),
    .Z(resp_msg[11]));
 BUF_X1 output40 (.A(net40),
    .Z(resp_msg[12]));
 BUF_X1 output41 (.A(net41),
    .Z(resp_msg[13]));
 BUF_X1 output42 (.A(net42),
    .Z(resp_msg[14]));
 BUF_X4 output43 (.A(net43),
    .Z(resp_msg[15]));
 BUF_X1 output44 (.A(net44),
    .Z(resp_msg[1]));
 BUF_X1 output45 (.A(net45),
    .Z(resp_msg[2]));
 BUF_X1 output46 (.A(net46),
    .Z(resp_msg[3]));
 BUF_X1 output47 (.A(net47),
    .Z(resp_msg[4]));
 BUF_X1 output48 (.A(net48),
    .Z(resp_msg[5]));
 BUF_X1 output49 (.A(net49),
    .Z(resp_msg[6]));
 BUF_X1 output50 (.A(net50),
    .Z(resp_msg[7]));
 BUF_X1 output51 (.A(net51),
    .Z(resp_msg[8]));
 BUF_X1 output52 (.A(net52),
    .Z(resp_msg[9]));
 BUF_X1 output53 (.A(net53),
    .Z(resp_val));
 BUF_X4 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 BUF_X4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 BUF_X4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 BUF_X4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 CLKBUF_X1 rebuffer1 (.A(\dpath.a_lt_b$in0[6] ),
    .Z(net54));
 CLKBUF_X1 rebuffer2 (.A(\dpath.a_lt_b$in0[6] ),
    .Z(net55));
 CLKBUF_X1 rebuffer3 (.A(\dpath.a_lt_b$in0[6] ),
    .Z(net56));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X2 FILLER_0_57 ();
 FILLCELL_X16 FILLER_0_62 ();
 FILLCELL_X4 FILLER_0_78 ();
 FILLCELL_X1 FILLER_0_82 ();
 FILLCELL_X8 FILLER_0_86 ();
 FILLCELL_X1 FILLER_0_94 ();
 FILLCELL_X4 FILLER_0_98 ();
 FILLCELL_X8 FILLER_0_105 ();
 FILLCELL_X2 FILLER_0_113 ();
 FILLCELL_X1 FILLER_0_115 ();
 FILLCELL_X8 FILLER_0_119 ();
 FILLCELL_X4 FILLER_0_127 ();
 FILLCELL_X8 FILLER_0_134 ();
 FILLCELL_X4 FILLER_0_142 ();
 FILLCELL_X1 FILLER_0_146 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X2 FILLER_0_157 ();
 FILLCELL_X1 FILLER_0_159 ();
 FILLCELL_X16 FILLER_0_163 ();
 FILLCELL_X8 FILLER_0_179 ();
 FILLCELL_X2 FILLER_0_187 ();
 FILLCELL_X32 FILLER_0_192 ();
 FILLCELL_X32 FILLER_0_224 ();
 FILLCELL_X4 FILLER_0_256 ();
 FILLCELL_X2 FILLER_0_260 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_132 ();
 FILLCELL_X32 FILLER_1_164 ();
 FILLCELL_X32 FILLER_1_196 ();
 FILLCELL_X32 FILLER_1_228 ();
 FILLCELL_X2 FILLER_1_260 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X4 FILLER_2_257 ();
 FILLCELL_X1 FILLER_2_261 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_257 ();
 FILLCELL_X1 FILLER_3_261 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X1 FILLER_4_97 ();
 FILLCELL_X16 FILLER_4_101 ();
 FILLCELL_X16 FILLER_4_120 ();
 FILLCELL_X8 FILLER_4_136 ();
 FILLCELL_X4 FILLER_4_144 ();
 FILLCELL_X32 FILLER_4_151 ();
 FILLCELL_X32 FILLER_4_183 ();
 FILLCELL_X32 FILLER_4_215 ();
 FILLCELL_X8 FILLER_4_247 ();
 FILLCELL_X4 FILLER_4_255 ();
 FILLCELL_X2 FILLER_4_259 ();
 FILLCELL_X1 FILLER_4_261 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_49 ();
 FILLCELL_X1 FILLER_5_57 ();
 FILLCELL_X8 FILLER_5_61 ();
 FILLCELL_X4 FILLER_5_69 ();
 FILLCELL_X1 FILLER_5_73 ();
 FILLCELL_X4 FILLER_5_77 ();
 FILLCELL_X8 FILLER_5_84 ();
 FILLCELL_X16 FILLER_5_96 ();
 FILLCELL_X2 FILLER_5_112 ();
 FILLCELL_X1 FILLER_5_114 ();
 FILLCELL_X16 FILLER_5_122 ();
 FILLCELL_X8 FILLER_5_138 ();
 FILLCELL_X2 FILLER_5_146 ();
 FILLCELL_X32 FILLER_5_152 ();
 FILLCELL_X32 FILLER_5_184 ();
 FILLCELL_X32 FILLER_5_216 ();
 FILLCELL_X8 FILLER_5_248 ();
 FILLCELL_X4 FILLER_5_256 ();
 FILLCELL_X2 FILLER_5_260 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_49 ();
 FILLCELL_X1 FILLER_6_57 ();
 FILLCELL_X1 FILLER_6_84 ();
 FILLCELL_X4 FILLER_6_102 ();
 FILLCELL_X2 FILLER_6_106 ();
 FILLCELL_X1 FILLER_6_108 ();
 FILLCELL_X4 FILLER_6_135 ();
 FILLCELL_X2 FILLER_6_139 ();
 FILLCELL_X1 FILLER_6_141 ();
 FILLCELL_X16 FILLER_6_166 ();
 FILLCELL_X4 FILLER_6_182 ();
 FILLCELL_X2 FILLER_6_186 ();
 FILLCELL_X1 FILLER_6_188 ();
 FILLCELL_X32 FILLER_6_197 ();
 FILLCELL_X32 FILLER_6_229 ();
 FILLCELL_X1 FILLER_6_261 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X2 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_74 ();
 FILLCELL_X2 FILLER_7_78 ();
 FILLCELL_X1 FILLER_7_80 ();
 FILLCELL_X4 FILLER_7_84 ();
 FILLCELL_X2 FILLER_7_88 ();
 FILLCELL_X1 FILLER_7_90 ();
 FILLCELL_X32 FILLER_7_96 ();
 FILLCELL_X16 FILLER_7_133 ();
 FILLCELL_X8 FILLER_7_152 ();
 FILLCELL_X2 FILLER_7_160 ();
 FILLCELL_X16 FILLER_7_165 ();
 FILLCELL_X4 FILLER_7_181 ();
 FILLCELL_X2 FILLER_7_185 ();
 FILLCELL_X8 FILLER_7_206 ();
 FILLCELL_X1 FILLER_7_214 ();
 FILLCELL_X8 FILLER_7_222 ();
 FILLCELL_X2 FILLER_7_230 ();
 FILLCELL_X1 FILLER_7_232 ();
 FILLCELL_X16 FILLER_7_236 ();
 FILLCELL_X8 FILLER_7_252 ();
 FILLCELL_X2 FILLER_7_260 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_60 ();
 FILLCELL_X2 FILLER_8_76 ();
 FILLCELL_X1 FILLER_8_78 ();
 FILLCELL_X4 FILLER_8_82 ();
 FILLCELL_X2 FILLER_8_86 ();
 FILLCELL_X16 FILLER_8_96 ();
 FILLCELL_X4 FILLER_8_112 ();
 FILLCELL_X1 FILLER_8_116 ();
 FILLCELL_X1 FILLER_8_127 ();
 FILLCELL_X8 FILLER_8_133 ();
 FILLCELL_X4 FILLER_8_141 ();
 FILLCELL_X2 FILLER_8_145 ();
 FILLCELL_X1 FILLER_8_147 ();
 FILLCELL_X8 FILLER_8_180 ();
 FILLCELL_X1 FILLER_8_188 ();
 FILLCELL_X1 FILLER_8_192 ();
 FILLCELL_X2 FILLER_8_196 ();
 FILLCELL_X8 FILLER_8_201 ();
 FILLCELL_X2 FILLER_8_209 ();
 FILLCELL_X1 FILLER_8_211 ();
 FILLCELL_X32 FILLER_8_229 ();
 FILLCELL_X1 FILLER_8_261 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_33 ();
 FILLCELL_X2 FILLER_9_41 ();
 FILLCELL_X1 FILLER_9_60 ();
 FILLCELL_X16 FILLER_9_63 ();
 FILLCELL_X1 FILLER_9_79 ();
 FILLCELL_X16 FILLER_9_94 ();
 FILLCELL_X1 FILLER_9_120 ();
 FILLCELL_X8 FILLER_9_138 ();
 FILLCELL_X4 FILLER_9_146 ();
 FILLCELL_X8 FILLER_9_160 ();
 FILLCELL_X4 FILLER_9_168 ();
 FILLCELL_X1 FILLER_9_172 ();
 FILLCELL_X8 FILLER_9_178 ();
 FILLCELL_X4 FILLER_9_186 ();
 FILLCELL_X2 FILLER_9_190 ();
 FILLCELL_X1 FILLER_9_196 ();
 FILLCELL_X2 FILLER_9_200 ();
 FILLCELL_X2 FILLER_9_212 ();
 FILLCELL_X2 FILLER_9_218 ();
 FILLCELL_X32 FILLER_9_226 ();
 FILLCELL_X4 FILLER_9_258 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_5 ();
 FILLCELL_X16 FILLER_10_9 ();
 FILLCELL_X4 FILLER_10_25 ();
 FILLCELL_X2 FILLER_10_42 ();
 FILLCELL_X2 FILLER_10_54 ();
 FILLCELL_X4 FILLER_10_64 ();
 FILLCELL_X1 FILLER_10_68 ();
 FILLCELL_X16 FILLER_10_87 ();
 FILLCELL_X4 FILLER_10_103 ();
 FILLCELL_X32 FILLER_10_124 ();
 FILLCELL_X32 FILLER_10_156 ();
 FILLCELL_X8 FILLER_10_188 ();
 FILLCELL_X4 FILLER_10_196 ();
 FILLCELL_X2 FILLER_10_200 ();
 FILLCELL_X32 FILLER_10_217 ();
 FILLCELL_X4 FILLER_10_249 ();
 FILLCELL_X2 FILLER_10_253 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_33 ();
 FILLCELL_X1 FILLER_11_35 ();
 FILLCELL_X16 FILLER_11_53 ();
 FILLCELL_X4 FILLER_11_69 ();
 FILLCELL_X2 FILLER_11_73 ();
 FILLCELL_X4 FILLER_11_77 ();
 FILLCELL_X2 FILLER_11_81 ();
 FILLCELL_X1 FILLER_11_83 ();
 FILLCELL_X32 FILLER_11_87 ();
 FILLCELL_X32 FILLER_11_119 ();
 FILLCELL_X32 FILLER_11_151 ();
 FILLCELL_X8 FILLER_11_183 ();
 FILLCELL_X4 FILLER_11_191 ();
 FILLCELL_X2 FILLER_11_195 ();
 FILLCELL_X1 FILLER_11_197 ();
 FILLCELL_X2 FILLER_11_202 ();
 FILLCELL_X1 FILLER_11_211 ();
 FILLCELL_X8 FILLER_11_221 ();
 FILLCELL_X2 FILLER_11_232 ();
 FILLCELL_X1 FILLER_11_241 ();
 FILLCELL_X2 FILLER_11_259 ();
 FILLCELL_X1 FILLER_11_261 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_49 ();
 FILLCELL_X1 FILLER_12_57 ();
 FILLCELL_X8 FILLER_12_65 ();
 FILLCELL_X4 FILLER_12_73 ();
 FILLCELL_X32 FILLER_12_82 ();
 FILLCELL_X32 FILLER_12_114 ();
 FILLCELL_X8 FILLER_12_146 ();
 FILLCELL_X2 FILLER_12_154 ();
 FILLCELL_X1 FILLER_12_163 ();
 FILLCELL_X16 FILLER_12_175 ();
 FILLCELL_X4 FILLER_12_191 ();
 FILLCELL_X1 FILLER_12_195 ();
 FILLCELL_X1 FILLER_12_242 ();
 FILLCELL_X1 FILLER_12_252 ();
 FILLCELL_X4 FILLER_12_256 ();
 FILLCELL_X2 FILLER_12_260 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X2 FILLER_13_13 ();
 FILLCELL_X1 FILLER_13_15 ();
 FILLCELL_X4 FILLER_13_19 ();
 FILLCELL_X2 FILLER_13_23 ();
 FILLCELL_X1 FILLER_13_35 ();
 FILLCELL_X1 FILLER_13_57 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_117 ();
 FILLCELL_X16 FILLER_13_127 ();
 FILLCELL_X8 FILLER_13_143 ();
 FILLCELL_X1 FILLER_13_151 ();
 FILLCELL_X16 FILLER_13_171 ();
 FILLCELL_X8 FILLER_13_187 ();
 FILLCELL_X4 FILLER_13_195 ();
 FILLCELL_X2 FILLER_13_199 ();
 FILLCELL_X16 FILLER_13_218 ();
 FILLCELL_X8 FILLER_13_238 ();
 FILLCELL_X4 FILLER_13_255 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X8 FILLER_14_14 ();
 FILLCELL_X2 FILLER_14_22 ();
 FILLCELL_X2 FILLER_14_27 ();
 FILLCELL_X1 FILLER_14_46 ();
 FILLCELL_X32 FILLER_14_66 ();
 FILLCELL_X32 FILLER_14_98 ();
 FILLCELL_X16 FILLER_14_130 ();
 FILLCELL_X8 FILLER_14_146 ();
 FILLCELL_X4 FILLER_14_154 ();
 FILLCELL_X2 FILLER_14_158 ();
 FILLCELL_X1 FILLER_14_160 ();
 FILLCELL_X8 FILLER_14_164 ();
 FILLCELL_X1 FILLER_14_172 ();
 FILLCELL_X1 FILLER_14_177 ();
 FILLCELL_X8 FILLER_14_181 ();
 FILLCELL_X32 FILLER_14_192 ();
 FILLCELL_X32 FILLER_14_224 ();
 FILLCELL_X4 FILLER_14_256 ();
 FILLCELL_X2 FILLER_14_260 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_21 ();
 FILLCELL_X32 FILLER_15_41 ();
 FILLCELL_X32 FILLER_15_73 ();
 FILLCELL_X32 FILLER_15_105 ();
 FILLCELL_X16 FILLER_15_137 ();
 FILLCELL_X8 FILLER_15_153 ();
 FILLCELL_X2 FILLER_15_161 ();
 FILLCELL_X1 FILLER_15_163 ();
 FILLCELL_X8 FILLER_15_181 ();
 FILLCELL_X4 FILLER_15_189 ();
 FILLCELL_X2 FILLER_15_203 ();
 FILLCELL_X8 FILLER_15_217 ();
 FILLCELL_X1 FILLER_15_225 ();
 FILLCELL_X2 FILLER_15_248 ();
 FILLCELL_X1 FILLER_15_250 ();
 FILLCELL_X4 FILLER_15_254 ();
 FILLCELL_X1 FILLER_15_258 ();
 FILLCELL_X2 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_6 ();
 FILLCELL_X1 FILLER_16_8 ();
 FILLCELL_X8 FILLER_16_15 ();
 FILLCELL_X4 FILLER_16_23 ();
 FILLCELL_X8 FILLER_16_34 ();
 FILLCELL_X1 FILLER_16_46 ();
 FILLCELL_X2 FILLER_16_50 ();
 FILLCELL_X32 FILLER_16_58 ();
 FILLCELL_X8 FILLER_16_90 ();
 FILLCELL_X2 FILLER_16_98 ();
 FILLCELL_X1 FILLER_16_100 ();
 FILLCELL_X32 FILLER_16_108 ();
 FILLCELL_X16 FILLER_16_140 ();
 FILLCELL_X8 FILLER_16_156 ();
 FILLCELL_X1 FILLER_16_164 ();
 FILLCELL_X8 FILLER_16_175 ();
 FILLCELL_X4 FILLER_16_183 ();
 FILLCELL_X2 FILLER_16_187 ();
 FILLCELL_X1 FILLER_16_198 ();
 FILLCELL_X1 FILLER_16_202 ();
 FILLCELL_X1 FILLER_16_206 ();
 FILLCELL_X2 FILLER_16_216 ();
 FILLCELL_X2 FILLER_16_223 ();
 FILLCELL_X1 FILLER_16_225 ();
 FILLCELL_X4 FILLER_16_229 ();
 FILLCELL_X2 FILLER_16_233 ();
 FILLCELL_X1 FILLER_16_235 ();
 FILLCELL_X2 FILLER_16_243 ();
 FILLCELL_X8 FILLER_16_248 ();
 FILLCELL_X4 FILLER_16_256 ();
 FILLCELL_X2 FILLER_16_260 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X8 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_17 ();
 FILLCELL_X1 FILLER_17_44 ();
 FILLCELL_X16 FILLER_17_68 ();
 FILLCELL_X8 FILLER_17_84 ();
 FILLCELL_X4 FILLER_17_92 ();
 FILLCELL_X2 FILLER_17_96 ();
 FILLCELL_X32 FILLER_17_117 ();
 FILLCELL_X4 FILLER_17_149 ();
 FILLCELL_X1 FILLER_17_153 ();
 FILLCELL_X16 FILLER_17_178 ();
 FILLCELL_X4 FILLER_17_194 ();
 FILLCELL_X2 FILLER_17_198 ();
 FILLCELL_X1 FILLER_17_200 ();
 FILLCELL_X4 FILLER_17_206 ();
 FILLCELL_X2 FILLER_17_210 ();
 FILLCELL_X2 FILLER_17_218 ();
 FILLCELL_X8 FILLER_17_230 ();
 FILLCELL_X1 FILLER_17_238 ();
 FILLCELL_X1 FILLER_17_246 ();
 FILLCELL_X2 FILLER_17_249 ();
 FILLCELL_X1 FILLER_17_251 ();
 FILLCELL_X1 FILLER_17_255 ();
 FILLCELL_X2 FILLER_17_259 ();
 FILLCELL_X1 FILLER_17_261 ();
 FILLCELL_X1 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_5 ();
 FILLCELL_X4 FILLER_18_13 ();
 FILLCELL_X1 FILLER_18_17 ();
 FILLCELL_X1 FILLER_18_21 ();
 FILLCELL_X2 FILLER_18_26 ();
 FILLCELL_X1 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X1 FILLER_18_35 ();
 FILLCELL_X8 FILLER_18_39 ();
 FILLCELL_X4 FILLER_18_47 ();
 FILLCELL_X2 FILLER_18_51 ();
 FILLCELL_X4 FILLER_18_59 ();
 FILLCELL_X2 FILLER_18_63 ();
 FILLCELL_X1 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_84 ();
 FILLCELL_X16 FILLER_18_116 ();
 FILLCELL_X8 FILLER_18_132 ();
 FILLCELL_X16 FILLER_18_147 ();
 FILLCELL_X8 FILLER_18_163 ();
 FILLCELL_X2 FILLER_18_171 ();
 FILLCELL_X32 FILLER_18_177 ();
 FILLCELL_X8 FILLER_18_209 ();
 FILLCELL_X4 FILLER_18_217 ();
 FILLCELL_X2 FILLER_18_221 ();
 FILLCELL_X1 FILLER_18_223 ();
 FILLCELL_X1 FILLER_18_243 ();
 FILLCELL_X8 FILLER_18_247 ();
 FILLCELL_X4 FILLER_18_255 ();
 FILLCELL_X2 FILLER_18_259 ();
 FILLCELL_X1 FILLER_18_261 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_9 ();
 FILLCELL_X8 FILLER_19_13 ();
 FILLCELL_X8 FILLER_19_41 ();
 FILLCELL_X4 FILLER_19_49 ();
 FILLCELL_X2 FILLER_19_53 ();
 FILLCELL_X2 FILLER_19_66 ();
 FILLCELL_X16 FILLER_19_77 ();
 FILLCELL_X8 FILLER_19_93 ();
 FILLCELL_X1 FILLER_19_101 ();
 FILLCELL_X32 FILLER_19_105 ();
 FILLCELL_X32 FILLER_19_137 ();
 FILLCELL_X16 FILLER_19_169 ();
 FILLCELL_X2 FILLER_19_185 ();
 FILLCELL_X16 FILLER_19_191 ();
 FILLCELL_X4 FILLER_19_207 ();
 FILLCELL_X1 FILLER_19_211 ();
 FILLCELL_X8 FILLER_19_216 ();
 FILLCELL_X2 FILLER_19_224 ();
 FILLCELL_X1 FILLER_19_226 ();
 FILLCELL_X16 FILLER_19_231 ();
 FILLCELL_X8 FILLER_19_247 ();
 FILLCELL_X4 FILLER_19_255 ();
 FILLCELL_X2 FILLER_19_259 ();
 FILLCELL_X1 FILLER_19_261 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_65 ();
 FILLCELL_X2 FILLER_20_72 ();
 FILLCELL_X1 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_88 ();
 FILLCELL_X8 FILLER_20_96 ();
 FILLCELL_X1 FILLER_20_104 ();
 FILLCELL_X1 FILLER_20_107 ();
 FILLCELL_X2 FILLER_20_110 ();
 FILLCELL_X16 FILLER_20_125 ();
 FILLCELL_X4 FILLER_20_141 ();
 FILLCELL_X1 FILLER_20_145 ();
 FILLCELL_X16 FILLER_20_149 ();
 FILLCELL_X4 FILLER_20_165 ();
 FILLCELL_X2 FILLER_20_169 ();
 FILLCELL_X1 FILLER_20_171 ();
 FILLCELL_X4 FILLER_20_175 ();
 FILLCELL_X2 FILLER_20_179 ();
 FILLCELL_X1 FILLER_20_181 ();
 FILLCELL_X1 FILLER_20_184 ();
 FILLCELL_X2 FILLER_20_187 ();
 FILLCELL_X8 FILLER_20_198 ();
 FILLCELL_X4 FILLER_20_206 ();
 FILLCELL_X1 FILLER_20_210 ();
 FILLCELL_X16 FILLER_20_214 ();
 FILLCELL_X8 FILLER_20_230 ();
 FILLCELL_X16 FILLER_20_242 ();
 FILLCELL_X4 FILLER_20_258 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_21 ();
 FILLCELL_X4 FILLER_21_40 ();
 FILLCELL_X1 FILLER_21_44 ();
 FILLCELL_X1 FILLER_21_48 ();
 FILLCELL_X1 FILLER_21_55 ();
 FILLCELL_X4 FILLER_21_59 ();
 FILLCELL_X2 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_75 ();
 FILLCELL_X2 FILLER_21_83 ();
 FILLCELL_X2 FILLER_21_110 ();
 FILLCELL_X2 FILLER_21_115 ();
 FILLCELL_X1 FILLER_21_123 ();
 FILLCELL_X2 FILLER_21_128 ();
 FILLCELL_X2 FILLER_21_134 ();
 FILLCELL_X16 FILLER_21_139 ();
 FILLCELL_X8 FILLER_21_155 ();
 FILLCELL_X2 FILLER_21_163 ();
 FILLCELL_X1 FILLER_21_165 ();
 FILLCELL_X4 FILLER_21_201 ();
 FILLCELL_X2 FILLER_21_226 ();
 FILLCELL_X1 FILLER_21_228 ();
 FILLCELL_X4 FILLER_21_232 ();
 FILLCELL_X2 FILLER_21_236 ();
 FILLCELL_X1 FILLER_21_249 ();
 FILLCELL_X2 FILLER_21_253 ();
 FILLCELL_X1 FILLER_21_255 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X2 FILLER_22_13 ();
 FILLCELL_X2 FILLER_22_18 ();
 FILLCELL_X4 FILLER_22_31 ();
 FILLCELL_X2 FILLER_22_35 ();
 FILLCELL_X1 FILLER_22_52 ();
 FILLCELL_X16 FILLER_22_72 ();
 FILLCELL_X1 FILLER_22_88 ();
 FILLCELL_X16 FILLER_22_94 ();
 FILLCELL_X8 FILLER_22_110 ();
 FILLCELL_X4 FILLER_22_118 ();
 FILLCELL_X32 FILLER_22_128 ();
 FILLCELL_X1 FILLER_22_160 ();
 FILLCELL_X2 FILLER_22_178 ();
 FILLCELL_X1 FILLER_22_180 ();
 FILLCELL_X16 FILLER_22_184 ();
 FILLCELL_X4 FILLER_22_200 ();
 FILLCELL_X2 FILLER_22_204 ();
 FILLCELL_X2 FILLER_22_215 ();
 FILLCELL_X1 FILLER_22_217 ();
 FILLCELL_X2 FILLER_22_221 ();
 FILLCELL_X1 FILLER_22_226 ();
 FILLCELL_X8 FILLER_22_250 ();
 FILLCELL_X4 FILLER_22_258 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_5 ();
 FILLCELL_X4 FILLER_23_13 ();
 FILLCELL_X2 FILLER_23_17 ();
 FILLCELL_X4 FILLER_23_21 ();
 FILLCELL_X1 FILLER_23_25 ();
 FILLCELL_X8 FILLER_23_29 ();
 FILLCELL_X4 FILLER_23_37 ();
 FILLCELL_X16 FILLER_23_46 ();
 FILLCELL_X1 FILLER_23_65 ();
 FILLCELL_X4 FILLER_23_69 ();
 FILLCELL_X32 FILLER_23_79 ();
 FILLCELL_X4 FILLER_23_111 ();
 FILLCELL_X1 FILLER_23_115 ();
 FILLCELL_X16 FILLER_23_125 ();
 FILLCELL_X8 FILLER_23_141 ();
 FILLCELL_X4 FILLER_23_149 ();
 FILLCELL_X8 FILLER_23_174 ();
 FILLCELL_X1 FILLER_23_182 ();
 FILLCELL_X4 FILLER_23_200 ();
 FILLCELL_X16 FILLER_23_207 ();
 FILLCELL_X8 FILLER_23_223 ();
 FILLCELL_X4 FILLER_23_231 ();
 FILLCELL_X1 FILLER_23_235 ();
 FILLCELL_X4 FILLER_23_256 ();
 FILLCELL_X2 FILLER_23_260 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_33 ();
 FILLCELL_X1 FILLER_24_37 ();
 FILLCELL_X16 FILLER_24_41 ();
 FILLCELL_X4 FILLER_24_57 ();
 FILLCELL_X2 FILLER_24_61 ();
 FILLCELL_X1 FILLER_24_63 ();
 FILLCELL_X8 FILLER_24_68 ();
 FILLCELL_X4 FILLER_24_76 ();
 FILLCELL_X1 FILLER_24_80 ();
 FILLCELL_X2 FILLER_24_85 ();
 FILLCELL_X1 FILLER_24_87 ();
 FILLCELL_X8 FILLER_24_90 ();
 FILLCELL_X2 FILLER_24_98 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_145 ();
 FILLCELL_X4 FILLER_24_153 ();
 FILLCELL_X1 FILLER_24_157 ();
 FILLCELL_X8 FILLER_24_176 ();
 FILLCELL_X2 FILLER_24_184 ();
 FILLCELL_X1 FILLER_24_186 ();
 FILLCELL_X32 FILLER_24_192 ();
 FILLCELL_X32 FILLER_24_224 ();
 FILLCELL_X4 FILLER_24_256 ();
 FILLCELL_X2 FILLER_24_260 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_9 ();
 FILLCELL_X4 FILLER_25_13 ();
 FILLCELL_X2 FILLER_25_20 ();
 FILLCELL_X1 FILLER_25_22 ();
 FILLCELL_X8 FILLER_25_49 ();
 FILLCELL_X4 FILLER_25_57 ();
 FILLCELL_X1 FILLER_25_61 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_73 ();
 FILLCELL_X1 FILLER_25_75 ();
 FILLCELL_X8 FILLER_25_93 ();
 FILLCELL_X4 FILLER_25_101 ();
 FILLCELL_X1 FILLER_25_105 ();
 FILLCELL_X4 FILLER_25_110 ();
 FILLCELL_X2 FILLER_25_114 ();
 FILLCELL_X1 FILLER_25_116 ();
 FILLCELL_X2 FILLER_25_120 ();
 FILLCELL_X32 FILLER_25_124 ();
 FILLCELL_X1 FILLER_25_156 ();
 FILLCELL_X16 FILLER_25_166 ();
 FILLCELL_X2 FILLER_25_182 ();
 FILLCELL_X1 FILLER_25_184 ();
 FILLCELL_X16 FILLER_25_190 ();
 FILLCELL_X4 FILLER_25_206 ();
 FILLCELL_X2 FILLER_25_210 ();
 FILLCELL_X32 FILLER_25_229 ();
 FILLCELL_X1 FILLER_25_261 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_33 ();
 FILLCELL_X4 FILLER_26_41 ();
 FILLCELL_X2 FILLER_26_45 ();
 FILLCELL_X1 FILLER_26_47 ();
 FILLCELL_X8 FILLER_26_51 ();
 FILLCELL_X2 FILLER_26_59 ();
 FILLCELL_X1 FILLER_26_65 ();
 FILLCELL_X8 FILLER_26_69 ();
 FILLCELL_X4 FILLER_26_77 ();
 FILLCELL_X2 FILLER_26_81 ();
 FILLCELL_X16 FILLER_26_86 ();
 FILLCELL_X4 FILLER_26_102 ();
 FILLCELL_X2 FILLER_26_106 ();
 FILLCELL_X1 FILLER_26_108 ();
 FILLCELL_X16 FILLER_26_119 ();
 FILLCELL_X8 FILLER_26_135 ();
 FILLCELL_X16 FILLER_26_164 ();
 FILLCELL_X4 FILLER_26_180 ();
 FILLCELL_X2 FILLER_26_184 ();
 FILLCELL_X2 FILLER_26_190 ();
 FILLCELL_X1 FILLER_26_192 ();
 FILLCELL_X8 FILLER_26_196 ();
 FILLCELL_X4 FILLER_26_204 ();
 FILLCELL_X32 FILLER_26_228 ();
 FILLCELL_X2 FILLER_26_260 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X16 FILLER_27_33 ();
 FILLCELL_X4 FILLER_27_49 ();
 FILLCELL_X2 FILLER_27_53 ();
 FILLCELL_X4 FILLER_27_72 ();
 FILLCELL_X1 FILLER_27_76 ();
 FILLCELL_X16 FILLER_27_84 ();
 FILLCELL_X4 FILLER_27_100 ();
 FILLCELL_X2 FILLER_27_104 ();
 FILLCELL_X1 FILLER_27_106 ();
 FILLCELL_X16 FILLER_27_129 ();
 FILLCELL_X2 FILLER_27_145 ();
 FILLCELL_X16 FILLER_27_149 ();
 FILLCELL_X8 FILLER_27_165 ();
 FILLCELL_X4 FILLER_27_173 ();
 FILLCELL_X2 FILLER_27_177 ();
 FILLCELL_X32 FILLER_27_196 ();
 FILLCELL_X32 FILLER_27_228 ();
 FILLCELL_X2 FILLER_27_260 ();
 FILLCELL_X2 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_3 ();
 FILLCELL_X32 FILLER_28_7 ();
 FILLCELL_X16 FILLER_28_39 ();
 FILLCELL_X4 FILLER_28_55 ();
 FILLCELL_X2 FILLER_28_59 ();
 FILLCELL_X1 FILLER_28_61 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X16 FILLER_28_97 ();
 FILLCELL_X1 FILLER_28_113 ();
 FILLCELL_X16 FILLER_28_118 ();
 FILLCELL_X8 FILLER_28_134 ();
 FILLCELL_X2 FILLER_28_142 ();
 FILLCELL_X1 FILLER_28_144 ();
 FILLCELL_X1 FILLER_28_154 ();
 FILLCELL_X16 FILLER_28_157 ();
 FILLCELL_X8 FILLER_28_173 ();
 FILLCELL_X4 FILLER_28_181 ();
 FILLCELL_X1 FILLER_28_185 ();
 FILLCELL_X32 FILLER_28_189 ();
 FILLCELL_X32 FILLER_28_221 ();
 FILLCELL_X8 FILLER_28_253 ();
 FILLCELL_X1 FILLER_28_261 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_97 ();
 FILLCELL_X1 FILLER_29_113 ();
 FILLCELL_X8 FILLER_29_117 ();
 FILLCELL_X2 FILLER_29_125 ();
 FILLCELL_X1 FILLER_29_127 ();
 FILLCELL_X1 FILLER_29_156 ();
 FILLCELL_X32 FILLER_29_176 ();
 FILLCELL_X32 FILLER_29_208 ();
 FILLCELL_X16 FILLER_29_240 ();
 FILLCELL_X4 FILLER_29_256 ();
 FILLCELL_X2 FILLER_29_260 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X16 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_153 ();
 FILLCELL_X32 FILLER_30_185 ();
 FILLCELL_X32 FILLER_30_217 ();
 FILLCELL_X8 FILLER_30_249 ();
 FILLCELL_X4 FILLER_30_257 ();
 FILLCELL_X1 FILLER_30_261 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X4 FILLER_31_257 ();
 FILLCELL_X1 FILLER_31_261 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X8 FILLER_32_129 ();
 FILLCELL_X4 FILLER_32_137 ();
 FILLCELL_X2 FILLER_32_141 ();
 FILLCELL_X1 FILLER_32_143 ();
 FILLCELL_X32 FILLER_32_148 ();
 FILLCELL_X32 FILLER_32_180 ();
 FILLCELL_X32 FILLER_32_212 ();
 FILLCELL_X16 FILLER_32_244 ();
 FILLCELL_X2 FILLER_32_260 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_97 ();
 FILLCELL_X8 FILLER_33_113 ();
 FILLCELL_X2 FILLER_33_121 ();
 FILLCELL_X16 FILLER_33_126 ();
 FILLCELL_X4 FILLER_33_142 ();
 FILLCELL_X32 FILLER_33_149 ();
 FILLCELL_X4 FILLER_33_181 ();
 FILLCELL_X1 FILLER_33_185 ();
 FILLCELL_X32 FILLER_33_189 ();
 FILLCELL_X32 FILLER_33_221 ();
 FILLCELL_X8 FILLER_33_253 ();
 FILLCELL_X1 FILLER_33_261 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_33 ();
 FILLCELL_X8 FILLER_34_49 ();
 FILLCELL_X4 FILLER_34_57 ();
 FILLCELL_X2 FILLER_34_61 ();
 FILLCELL_X8 FILLER_34_66 ();
 FILLCELL_X4 FILLER_34_74 ();
 FILLCELL_X2 FILLER_34_78 ();
 FILLCELL_X1 FILLER_34_80 ();
 FILLCELL_X16 FILLER_34_84 ();
 FILLCELL_X8 FILLER_34_100 ();
 FILLCELL_X4 FILLER_34_108 ();
 FILLCELL_X2 FILLER_34_118 ();
 FILLCELL_X1 FILLER_34_120 ();
 FILLCELL_X16 FILLER_34_124 ();
 FILLCELL_X2 FILLER_34_140 ();
 FILLCELL_X2 FILLER_34_148 ();
 FILLCELL_X32 FILLER_34_153 ();
 FILLCELL_X1 FILLER_34_185 ();
 FILLCELL_X32 FILLER_34_189 ();
 FILLCELL_X32 FILLER_34_221 ();
 FILLCELL_X8 FILLER_34_253 ();
 FILLCELL_X1 FILLER_34_261 ();
endmodule
